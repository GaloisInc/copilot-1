package FloatsTypes where {
import FloatingPoint;
                    
import Vector
}