import FloatingPoint::*;

import "BDPI" function Float bs_fp_expf (Float x);
import "BDPI" function Double bs_fp_exp (Double x);
import "BDPI" function Float bs_fp_logf (Float x);
import "BDPI" function Double bs_fp_log (Double x);
import "BDPI" function Float bs_fp_acosf (Float x);
import "BDPI" function Double bs_fp_acos (Double x);
import "BDPI" function Float bs_fp_asinf (Float x);
import "BDPI" function Double bs_fp_asin (Double x);
import "BDPI" function Float bs_fp_atanf (Float x);
import "BDPI" function Double bs_fp_atan (Double x);
import "BDPI" function Float bs_fp_cosf (Float x);
import "BDPI" function Double bs_fp_cos (Double x);
import "BDPI" function Float bs_fp_sinf (Float x);
import "BDPI" function Double bs_fp_sin (Double x);
import "BDPI" function Float bs_fp_tanf (Float x);
import "BDPI" function Double bs_fp_tan (Double x);
import "BDPI" function Float bs_fp_acoshf (Float x);
import "BDPI" function Double bs_fp_acosh (Double x);
import "BDPI" function Float bs_fp_asinhf (Float x);
import "BDPI" function Double bs_fp_asinh (Double x);
import "BDPI" function Float bs_fp_atanhf (Float x);
import "BDPI" function Double bs_fp_atanh (Double x);
import "BDPI" function Float bs_fp_coshf (Float x);
import "BDPI" function Double bs_fp_cosh (Double x);
import "BDPI" function Float bs_fp_sinhf (Float x);
import "BDPI" function Double bs_fp_sinh (Double x);
import "BDPI" function Float bs_fp_tanhf (Float x);
import "BDPI" function Double bs_fp_tanh (Double x);
import "BDPI" function Float bs_fp_ceilf (Float x);
import "BDPI" function Double bs_fp_ceil (Double x);
import "BDPI" function Float bs_fp_floorf (Float x);
import "BDPI" function Double bs_fp_floor (Double x);
import "BDPI" function Float bs_fp_sqrtf (Float x);
import "BDPI" function Double bs_fp_sqrt (Double x);
import "BDPI" function Float bs_fp_powf (Float x, Float y);
import "BDPI" function Double bs_fp_pow (Double x, Double y);
import "BDPI" function Float bs_fp_atan2f (Float x, Float y);
import "BDPI" function Double bs_fp_atan2 (Double x, Double y);
import "BDPI" function Float bs_fp_logbf (Float x, Float y);
import "BDPI" function Double bs_fp_logb (Double x, Double y);
