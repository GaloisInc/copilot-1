package Floats where {
import FloatingPoint;
                    
import Vector;
             
import FloatsTypes;
                  
import BluespecFP;
                 
interface FloatsIfc {-# always_ready , always_enabled  #-} = {
    rtf_guard :: Prelude.Bool;
    rtf_arg0 :: Float;
    rtf_arg1 :: Float;
    rtf_arg2 :: Float
};
 
{-# properties mkFloats = { verilog } #-};
                                         
mkFloats :: Prelude.Module FloatsIfc;
mkFloats = 
    module {
      s0_0 :: Prelude.Reg Float <- mkReg (5.104235503814077e38::Float);
      let { s0 :: Vector.Vector 1 (Prelude.Reg Float);
            s0 =  update newVector 0 s0_0; };
      s1_0 :: Prelude.Reg Float <- mkReg (3.402823669209385e38::Float);
      s1_1 :: Prelude.Reg Float <- mkReg
                                     ((Prelude.negate 3.402823669209385e38)::Float);
      let { s1 :: Vector.Vector 2 (Prelude.Reg Float);
            s1 =  update (update newVector 0 s1_0) 1 s1_1; };
      s2_0 :: Prelude.Reg Float <- mkReg (0.0::Float);
      s2_1 :: Prelude.Reg Float <- mkReg (0.0::Float);
      let { s2 :: Vector.Vector 2 (Prelude.Reg Float);
            s2 =  update (update newVector 0 s2_0) 1 s2_1; };
      s0_idx :: Prelude.Reg (Prelude.Bit 64) <- mkReg 0;
      s1_idx :: Prelude.Reg (Prelude.Bit 64) <- mkReg 0;
      s2_idx :: Prelude.Reg (Prelude.Bit 64) <- mkReg 0;
      let { s0_get :: Prelude.Bit 64 -> Float;
            s0_get x =  (select s0 ((Prelude.%) ((+) s0_idx x) 1))._read;
            s1_get :: Prelude.Bit 64 -> Float;
            s1_get x =  (select s1 ((Prelude.%) ((+) s1_idx x) 2))._read;
            s2_get :: Prelude.Bit 64 -> Float;
            s2_get x =  (select s2 ((Prelude.%) ((+) s2_idx x) 2))._read;
            s0_gen :: Float;
            s0_gen =  s0_get 0;
            s1_gen :: Float;
            s1_gen =  s1_get 0;
            s2_gen :: Float;
            s2_gen =  s2_get 0; };
      rules {
        
        "step":  when Prelude.True
                  ==>
                    action { (select s0 s0_idx) := s0_gen;
                             (select s1 s1_idx) := s1_gen;
                             (select s2 s2_idx) := s2_gen;
                             s0_idx := (Prelude.%) ((+) s0_idx 1) 1;
                             s1_idx := (Prelude.%) ((+) s1_idx 1) 2;
                             s2_idx := (Prelude.%) ((+) s2_idx 1) 2;
                             }
      };
      Prelude.return
        (interface FloatsIfc {
           rtf_guard :: Prelude.Bool;
           rtf_guard =  Prelude.True;;
           rtf_arg0 :: Float;
           rtf_arg0 =  s0_get 0;;
           rtf_arg1 :: Float;
           rtf_arg1 =  s1_get 0;;
           rtf_arg2 :: Float;
           rtf_arg2 =  s2_get 0;
         })
    };;
      
interface FloatsRulesIfc = {
    rtf_action :: Float -> Float -> Float -> Prelude.Action
};
 
mkFloatsRules :: FloatsIfc -> FloatsRulesIfc -> Prelude.Rules;
mkFloatsRules ifc ifcRules = 
    rules {
      
      "rtf":  when ifc.rtf_guard
               ==>
                 ifcRules.rtf_action ifc.rtf_arg0 ifc.rtf_arg1 ifc.rtf_arg2
    };;
      
addFloatsRules :: FloatsIfc ->
                  FloatsRulesIfc -> Prelude.Module Prelude.Empty;
addFloatsRules ifc ifcRules = 
    Prelude.addRules (mkFloatsRules ifc ifcRules);
}